
module vprom(input clk,
	     input 	  reset,
	     input [7:0]  a,
	     output [3:0] d);

   reg [3:0] q;

   assign d = q;
   
   always @(posedge clk)
     case (a)
	8'h00: q = 4'b0000;
	8'h01: q = 4'b0000;
	8'h02: q = 4'b0000;
	8'h03: q = 4'b0000;
	8'h04: q = 4'b0000;
	8'h05: q = 4'b0000;
	8'h06: q = 4'b0000;
	8'h07: q = 4'b0000;
	8'h08: q = 4'b0000;
	8'h09: q = 4'b0000;
	8'h0a: q = 4'b0000;
	8'h0b: q = 4'b0000;
	8'h0c: q = 4'b0000;
	8'h0d: q = 4'b0000;
	8'h0e: q = 4'b0000;
	8'h0f: q = 4'b0000;
	8'h10: q = 4'b0000;
	8'h11: q = 4'b0000;
	8'h12: q = 4'b0000;
	8'h13: q = 4'b0000;
	8'h14: q = 4'b0000;
	8'h15: q = 4'b0000;
	8'h16: q = 4'b0000;
	8'h17: q = 4'b0000;
	8'h18: q = 4'b0000;
	8'h19: q = 4'b0000;
	8'h1a: q = 4'b0000;
	8'h1b: q = 4'b0000;
	8'h1c: q = 4'b0000;
	8'h1d: q = 4'b0000;
	8'h1e: q = 4'b0000;
	8'h1f: q = 4'b0000;
	8'h20: q = 4'b0000;
	8'h21: q = 4'b0000;
	8'h22: q = 4'b0000;
	8'h23: q = 4'b0000;
	8'h24: q = 4'b0000;
	8'h25: q = 4'b0000;
	8'h26: q = 4'b0000;
	8'h27: q = 4'b0000;
	8'h28: q = 4'b0000;
	8'h29: q = 4'b0000;
	8'h2a: q = 4'b0000;
	8'h2b: q = 4'b0000;
	8'h2c: q = 4'b0000;
	8'h2d: q = 4'b0000;
	8'h2e: q = 4'b0000;
	8'h2f: q = 4'b0000;
	8'h30: q = 4'b0000;
	8'h31: q = 4'b0000;
	8'h32: q = 4'b0000;
	8'h33: q = 4'b0000;
	8'h34: q = 4'b0000;
	8'h35: q = 4'b0000;
	8'h36: q = 4'b0000;
	8'h37: q = 4'b0000;
	8'h38: q = 4'b0000;
	8'h39: q = 4'b0000;
	8'h3a: q = 4'b0000;
	8'h3b: q = 4'b0000;
	8'h3c: q = 4'b0000;
	8'h3d: q = 4'b0000;
	8'h3e: q = 4'b0000;
	8'h3f: q = 4'b0000;
	8'h40: q = 4'b0000;
	8'h41: q = 4'b0000;
	8'h42: q = 4'b0000;
	8'h43: q = 4'b0000;
	8'h44: q = 4'b0000;
	8'h45: q = 4'b0000;
	8'h46: q = 4'b0000;
	8'h47: q = 4'b0000;
	8'h48: q = 4'b0000;
	8'h49: q = 4'b0000;
	8'h4a: q = 4'b0000;
	8'h4b: q = 4'b0000;
	8'h4c: q = 4'b0000;
	8'h4d: q = 4'b0000;
	8'h4e: q = 4'b0000;
	8'h4f: q = 4'b0000;
	8'h50: q = 4'b0000;
	8'h51: q = 4'b0000;
	8'h52: q = 4'b0000;
	8'h53: q = 4'b0000;
	8'h54: q = 4'b0000;
	8'h55: q = 4'b0000;
	8'h56: q = 4'b0000;
	8'h57: q = 4'b0000;
	8'h58: q = 4'b0000;
	8'h59: q = 4'b0000;
	8'h5a: q = 4'b0000;
	8'h5b: q = 4'b0000;
	8'h5c: q = 4'b0000;
	8'h5d: q = 4'b0000;
	8'h5e: q = 4'b0000;
	8'h5f: q = 4'b0000;
	8'h60: q = 4'b0000;
	8'h61: q = 4'b0000;
	8'h62: q = 4'b0000;
	8'h63: q = 4'b0000;
	8'h64: q = 4'b0000;
	8'h65: q = 4'b0000;
	8'h66: q = 4'b0000;
	8'h67: q = 4'b0000;
	8'h68: q = 4'b0010;
	8'h69: q = 4'b0010;
	8'h6a: q = 4'b0010;
	8'h6b: q = 4'b0010;
	8'h6c: q = 4'b0010;
	8'h6d: q = 4'b0010;
	8'h6e: q = 4'b0010;
	8'h6f: q = 4'b0010;
	8'h70: q = 4'b0010;
	8'h71: q = 4'b0010;
	8'h72: q = 4'b0010;
	8'h73: q = 4'b0010;
	8'h74: q = 4'b0010;
	8'h75: q = 4'b0010;
	8'h76: q = 4'b0010;
	8'h77: q = 4'b0010;
	8'h78: q = 4'b0010;
	8'h79: q = 4'b0010;
	8'h7a: q = 4'b0010;
	8'h7b: q = 4'b0010;
	8'h7c: q = 4'b0010;
	8'h7d: q = 4'b0010;
	8'h7e: q = 4'b0010;
	8'h7f: q = 4'b1010;
	8'h80: q = 4'b0000;
	8'h81: q = 4'b1010;
	8'h82: q = 4'b1010;
	8'h83: q = 4'b1010;
	8'h84: q = 4'b1010;
	8'h85: q = 4'b1110;
	8'h86: q = 4'b0000;
	8'h87: q = 4'b0000;
	8'h88: q = 4'b0000;
	8'h89: q = 4'b0000;
	8'h8a: q = 4'b0000;
	8'h8b: q = 4'b0000;
	8'h8c: q = 4'b0000;
	8'h8d: q = 4'b0000;
	8'h8e: q = 4'b0000;
	8'h8f: q = 4'b0000;
	8'h90: q = 4'b0000;
	8'h91: q = 4'b0000;
	8'h92: q = 4'b0000;
	8'h93: q = 4'b0000;
	8'h94: q = 4'b0000;
	8'h95: q = 4'b0000;
	8'h96: q = 4'b0000;
	8'h97: q = 4'b0000;
	8'h98: q = 4'b0000;
	8'h99: q = 4'b0000;
	8'h9a: q = 4'b0000;
	8'h9b: q = 4'b0000;
	8'h9c: q = 4'b0000;
	8'h9d: q = 4'b0000;
	8'h9e: q = 4'b0000;
	8'h9f: q = 4'b0000;
	8'ha0: q = 4'b0000;
	8'ha1: q = 4'b0000;
	8'ha2: q = 4'b0000;
	8'ha3: q = 4'b0000;
	8'ha4: q = 4'b0000;
	8'ha5: q = 4'b0000;
	8'ha6: q = 4'b0000;
	8'ha7: q = 4'b0000;
	8'ha8: q = 4'b0000;
	8'ha9: q = 4'b0000;
	8'haa: q = 4'b0000;
	8'hab: q = 4'b0000;
	8'hac: q = 4'b0000;
	8'had: q = 4'b0000;
	8'hae: q = 4'b0000;
	8'haf: q = 4'b0000;
	8'hb0: q = 4'b0000;
	8'hb1: q = 4'b0000;
	8'hb2: q = 4'b0000;
	8'hb3: q = 4'b0000;
	8'hb4: q = 4'b0000;
	8'hb5: q = 4'b0000;
	8'hb6: q = 4'b0000;
	8'hb7: q = 4'b0000;
	8'hb8: q = 4'b0000;
	8'hb9: q = 4'b0000;
	8'hba: q = 4'b0000;
	8'hbb: q = 4'b0000;
	8'hbc: q = 4'b0000;
	8'hbd: q = 4'b0000;
	8'hbe: q = 4'b0000;
	8'hbf: q = 4'b0000;
	8'hc0: q = 4'b0000;
	8'hc1: q = 4'b0000;
	8'hc2: q = 4'b0000;
	8'hc3: q = 4'b0000;
	8'hc4: q = 4'b0000;
	8'hc5: q = 4'b0000;
	8'hc6: q = 4'b0000;
	8'hc7: q = 4'b0000;
	8'hc8: q = 4'b0000;
	8'hc9: q = 4'b0000;
	8'hca: q = 4'b0000;
	8'hcb: q = 4'b0000;
	8'hcc: q = 4'b0000;
	8'hcd: q = 4'b0000;
	8'hce: q = 4'b0000;
	8'hcf: q = 4'b0000;
	8'hd0: q = 4'b0000;
	8'hd1: q = 4'b0000;
	8'hd2: q = 4'b0000;
	8'hd3: q = 4'b0000;
	8'hd4: q = 4'b0000;
	8'hd5: q = 4'b0000;
	8'hd6: q = 4'b0000;
	8'hd7: q = 4'b0000;
	8'hd8: q = 4'b0000;
	8'hd9: q = 4'b0000;
	8'hda: q = 4'b0000;
	8'hdb: q = 4'b0000;
	8'hdc: q = 4'b0000;
	8'hdd: q = 4'b0000;
	8'hde: q = 4'b0000;
	8'hdf: q = 4'b0000;
	8'he0: q = 4'b1010;
	8'he1: q = 4'b1010;
	8'he2: q = 4'b1010;
	8'he3: q = 4'b1010;
	8'he4: q = 4'b1010;
	8'he5: q = 4'b1010;
	8'he6: q = 4'b1010;
	8'he7: q = 4'b1010;
	8'he8: q = 4'b1010;
	8'he9: q = 4'b1010;
	8'hea: q = 4'b1010;
	8'heb: q = 4'b1010;
	8'hec: q = 4'b1010;
	8'hed: q = 4'b1010;
	8'hee: q = 4'b1010;
	8'hef: q = 4'b1010;
	8'hf0: q = 4'b1010;
	8'hf1: q = 4'b1010;
	8'hf2: q = 4'b1011;
	8'hf3: q = 4'b1011;
	8'hf4: q = 4'b1011;
	8'hf5: q = 4'b1010;
	8'hf6: q = 4'b1010;
	8'hf7: q = 4'b1010;
	8'hf8: q = 4'b1010;
	8'hf9: q = 4'b1010;
	8'hfa: q = 4'b1010;
	8'hfb: q = 4'b1010;
	8'hfc: q = 4'b1010;
	8'hfd: q = 4'b1010;
	8'hfe: q = 4'b1010;
	8'hff: q = 4'b1010;
     endcase
   
endmodule // vprom

